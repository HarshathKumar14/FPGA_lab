


module twobitmul(
input [1:0]a,b,

output [3:0]c
    );
    
    assign c=a*b;
endmodule
